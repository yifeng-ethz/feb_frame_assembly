alt_parallel_add_inst : alt_parallel_add PORT MAP (
		clock	 => clock_sig,
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		data2x	 => data2x_sig,
		data3x	 => data3x_sig,
		result	 => result_sig
	);
